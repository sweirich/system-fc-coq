Require Import Omega.

Require Export Typing.
Require Export Coq.Logic.Decidable.

Module WEAKENING.
Import SYSTEMFC.
Import SHIFTING.
Import SUBSTITUTION.
Import TYPING.

(** This module contains various properties related to 
    Weakening and Strengthening for the type system. 
  
*)


(* ####################################################### *)  

(* ####################################################### *)  
